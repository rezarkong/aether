library ieee;
use ieee.std_logic_1164.all;

package enae_pkg is

    type state0_t_arr is array (0 to 3) of std_logic_vector(127 downto 0);
    type state1_t_arr is array (0 to 5) of std_logic_vector(127 downto 0);
    type state2_t_arr is array (0 to 8) of std_logic_vector(127 downto 0);
   
end package;
